module ROM (
input logic [5:0] address, // 16 addresses in total
output logic [63:0] data); // 8bits/address
always_comb
begin  
case (address)
0:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		1:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		2:data=64'b1111111111111111111111111111111110111111111111111111111111111111;
		3:data=64'b1111111111111111111111111111111101011111111111111111111111111111;
		4:data=64'b1111111111111111111111111111111110111111111111111111111111111111;
		5:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		6:data=64'b1111111111111000000000001111111111111111000000000000111111111111;
		7:data=64'b1111111111100000000000000011111111111100000000000000001111111111;
		8:data=64'b1111111110000000000000000000111111110000000000000000000011111111;
		9:data=64'b1111111000000000000000000000011111100000000000000000000000111111;
		10:data=64'b1111000000000000000000000000001110000000000000000000000000001111;
		11:data=64'b1110000000000000000000000000000100000000000000000000000000000111;
		12:data=64'b1100000000000000000000000000000000000000000000000000000000000011;
		13:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		14:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		15:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		16:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		17:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		18:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		19:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		20:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		21:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		22:data=64'b1000000000000000000000000000000000000000000000000000000000000001;
		23:data=64'b1100000000000000000000000000000000000000000000000000000000000011;
		24:data=64'b1110000000000000000000000000000000000000000000000000000000000111;
		25:data=64'b1111000000000000000000000000000000000000000000000000000000001111;
		26:data=64'b1111110000000000000000000000000000000000000000000000000000111111;
		27:data=64'b1111111100000000000000000000000000000000000000000000000011111111;
		28:data=64'b1111111111000000000000000000000000000000000000000000001111111111;
		29:data=64'b1111111111110000000000000000000000000000000000000000111111111111;
		30:data=64'b1111111111111100000000000000000000000000000000000011111111111111;
		31:data=64'b1111111111111111000000000000000000000000000000001111111111111111;
		32:data=64'b1111111111111111110000000000000000000000000000111111111111111111;
		33:data=64'b1111111111111111111100000000000000000000000011111111111111111111;
		34:data=64'b1111111111111111111111000000000000000000001111111111111111111111;
		35:data=64'b1111111111111111111111110000000000000000111111111111111111111111;
		36:data=64'b1111111111111111111111111100000000000011111111111111111111111111;
		37:data=64'b1111111111111111111111111111100000001111111111111111111111111111;
		38:data=64'b1111111111111111111111111111111000111111111111111111111111111111;
		39:data=64'b1111111111111111111111111111111101111111111111111111111111111111;
		40:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		41:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		42:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		43:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		44:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		45:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		46:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		47:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		default:data=64'b1111111111111111111111111111111111111111111111111111111111111111;
		endcase
end
endmodule