module rom (
input logic [5:0] address, // 16 addresses in total
output logic [63:0] data); // 8bits/address
always_comb
begin  
case (address)
0 : data =64'b0000000000111100000000000110000000000000000000000000000001111100;
1 : data =64'b0000000000111100000000000000000001111100000000000000000000111100;
2 : data =64'b0000000000111100000001111100000000000000000000000000000000001100;
3 : data =64'b0000000001111100000000000000001111100000000000000000000000000111;
4 : data =64'b0000000001111100000000000000000000000000000000000000000000000111;
5 : data =64'b0000000000000000111111000000000000000000000000000000000000000111;
6 : data =64'b0000000000000000000001111110000000000000000000000000000000000111;
7 : data =64'b0000000000000000000001111110000000000000000000000000000000000111;
8 : data =64'b0000000000000000000001111110000000000000000000000000000000000111;
9 : data =64'b0000000000000000000001111110000000000000000000000000000000000111;
10 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
11 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
12 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
13 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
14: data =  64'b0000000000000000000111111000000000000000000000000000000000000111;
15 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
16 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
17 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
18 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
19 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
20 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
21 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
22 : data = 64'b0000000000000000000111111000000000000000000000000000000000000111;
23: data = 64'b1111111111111111111111100000111111111111111111111111111111111111;
24: data = 64'b1111111111111111111111100000111111111111111111111111111111111111;
25: data = 64'b1111111111111111111111100000111111111111111111111111111111111111;
26: data = 64'b1111111111111111111111100000111111111111111111111111111111111111;
27: data = 64'b1111111111111111111111100000111111111111111111111111111111111111;
28: data = 64'b1111111111111111111111100000111111111111111111111111111111111111;
29: data =  64'b0000000000000000000000000000000000000000000000000000000000000111;
30 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
31 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
32 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
33 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
34 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
35 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
36 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
37 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
38 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
39 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
40 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
41 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
42 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
43 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
44 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
45 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
46 : data = 64'b0000000000000000000000000000000000000000000000000000000000000111;
47 : data = 64'b0000000000000000000000000000000000000000000000000000000001111111;

default : data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
endcase;
end
endmodule