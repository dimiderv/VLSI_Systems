module rom (
input logic [5:0] address, // 16 addresses in total
output logic [63:0] data); // 8bits/address
always_comb
begin
case (address)
0 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
1 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
2 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
3 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
4 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
5 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
6 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
7 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
8 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
9 : data =64'b0001100000000000000011111000001111100001111110000011111000001111;
10 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
11 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
12 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
13 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
14: data =  64'b001100000000000000011111000001111100001111110000011111000001111;
15 : data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
16 : data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
17 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
18 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
19 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
20 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
21 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
22 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
23: data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
24: data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
25: data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
26: data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
27: data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
28: data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
29: data =  64'b0001100000000000000011111000001111100001111110000011111000001111;
30 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
31 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
32 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
33 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
34 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
35 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
36 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
37 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
38 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
39 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
40 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
41 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
42 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
43 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
44 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
45 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
46 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;
47 : data = 64'b0001100000000000000011111000001111100001111110000011111000001111;

default : data = 64'b1111111111111111111111111111111111111111111111111111111111111111;
endcase;
end
endmodule